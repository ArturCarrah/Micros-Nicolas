library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity control_unit is
    port (
        -- controle
        clk 
        rst
        we

        -- funcoes
        
    );
end entity;